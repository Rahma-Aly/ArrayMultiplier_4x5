`ifndef DEFINITIONS_SV
`define DEFINITIONS_SV


package definitions;
	parameter INPUT1_WIDTH = 4;

    parameter INPUT2_WIDTH = 5;

    
endpackage : definitions


`endif
